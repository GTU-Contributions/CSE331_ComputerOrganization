module bit32_alu_testbench();	
	reg  [3:0] ALUop;
	reg  [31:0]a;
	reg  [31:0]b;
	wire [31:0]r;
	wire Z, V, CarryOut;
	
	bit32_alu test(Z, V, CarryOut, r, a, b, ALUop);

initial begin

ALUop = 4'b0110; // A - B
a = 32'b00000000000000000000000000000010; // +2
b = 32'b00000000000000000000000000000001; // +1
#50;

ALUop = 4'b0110; // A - B
a = 32'b00000000000000000000000000000001; // +1
b = 32'b00000000000000000000000000000010; // +2
#50;

ALUop = 4'b0010; // A + B
a = 32'b00000000000000000000000000000101; // +5
b = 32'b00000000000000000000000000000110; // +6
#50;

ALUop = 4'b0110; // A - B
a = 32'b11111111111111111111111111111011; // -5
b = 32'b00000000000000000000000000000110; // +6
#50;

ALUop = 4'b0000; // A and B
a = 32'b01010101010101010101010101010101; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0000; // A and B
a = 32'b10101010101010101010101010101010; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0000; // A and B
a = 32'b11111111111111110000000000000000; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0001; // A or B
a = 32'b01010101010101010101010101010101; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0001; // A or B
a = 32'b10101010101010101010101010101010; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0001; // A or B
a = 32'b11111111111111110000000000000000; 
b = 32'b01000000000000000101010101010101;
#50;

ALUop = 4'b0010; // A + B
a = 32'b01010101010101010101010101010101; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0010; // A + B
a = 32'b10101010101010101010101010101010; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b0010; // A + B
a = 32'b10000000000000001111111111111111; 
b = 32'b11000000000000001010101010101010;
#50;

ALUop = 4'b1010; // A + B unsig
a = 32'b01010101010101010101010101010101; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b1010; // A + B unsig
a = 32'b10101010101010101010101010101010; 
b = 32'b01010101010101010101010101010101;
#50;

ALUop = 4'b1010; // A + B unsig
a = 32'b10000000000000001111111111111111; 
b = 32'b11000000000000001010101010101010;
#50;

ALUop = 4'b0110; // A - B
a = 32'b00000000000000001111111111111111; 
b = 32'b00000000000000001010101010101010;
#50;

ALUop = 4'b0110; // A - B
a = 32'b00000000000000001111111111111111; 
b = 32'b00000000000000011010101010101010;
#50;

ALUop = 4'b0110; // A - B
a = 32'b10000000000000001111111111111111; 
b = 32'b11000000000000001010101010101010;
#50;

ALUop = 4'b1110; // A - B unsig
a = 32'b00000000000000001111111111111111; 
b = 32'b00000000000000001010101010101010;
#50;

ALUop = 4'b1110; // A - B unsig
a = 32'b00000000000000001111111111111111; 
b = 32'b00000000000000011010101010101010;
#50;

ALUop = 4'b1110; // A - B unsig
a = 32'b10000000000000001111111111111111; 
b = 32'b11000000000000001010101010101010;
#50;

ALUop = 4'b0101; // A nor B
a = 32'b00000000000000011111111111111111; 
b = 32'b00000000000000000010101010101010;
#50;

ALUop = 4'b0101; // A nor B
a = 32'b00000000000000000010101010101010;
b = 32'b00000000000000011111111111111111;
#50;

ALUop = 4'b0111; // SLT
a = 32'b01111111111111111111111111111111; 
b = 32'b00000000000000000000000000000001;
#50;

ALUop = 4'b0111; // SLT
a = 32'b11111111111111111111111111111111; 
b = 32'b00000000000000000000000000000001;
#50;

ALUop = 4'b0111; // SLT
a = 32'b01000000000000000000010101010001; 
b = 32'b10000000111111111111111111111111;
#50;

ALUop = 4'b0111; // SLT
a = 32'b11000000000000000000000000000001; 
b = 32'b10000000000000000000000000000001;
#50;

ALUop = 4'b0111; // SLT
a = 32'b10010000000000000000000000000001; 
b = 32'b11000000000000000000000000000001;
#50;

ALUop = 4'b1111; // SLTU
a = 32'b01111111111111111111111111111111; 
b = 32'b00000000000000000000000000000001;
#50;

ALUop = 4'b1111; // SLTU
a = 32'b11111111111111111111111111111111; 
b = 32'b00000000000000000000000000000001;
#50;

ALUop = 4'b1111; // SLTU
a = 32'b01000000000000000000010101010001; 
b = 32'b10000000111111111111111111111111;
#50;

ALUop = 4'b1111; // SLTU
a = 32'b11000000000000000000000000000001; 
b = 32'b10000000000000000000000000000001;
#50;

ALUop = 4'b1111; // SLTU
a = 32'b10010000000000000000000000000001; 
b = 32'b11000000000000000000000000000001;
#50;

ALUop = 4'b1000; // SLL
a = 32'b01010101011111111111100001111100; 
b = 32'b00000000000000000000000000000001;
#50;

ALUop = 4'b1000; // SLL
a = 32'b01010100000000000000000010010011; 
b = 32'b10000000111111111111111111111111;
#50;

ALUop = 4'b1001; // SRL
a = 32'b11000000000000000000000001000001; 
b = 32'b10000000000000000000000000000001;
#50;

ALUop = 4'b1001; // SRL
a = 32'b10010000000000000000000010000001; 
b = 32'b11000000000000000000000000000001;
#50;

end
 
initial
begin
$monitor("ALUop=%4b,\n a=%32b,\n b=%32b,\n r=%32b,\n Z=%1b, V=%1b, C=%1b, ", ALUop, a, b, r, Z, V, CarryOut);
end
 
endmodule